module DontCareCase (
  output       out1,
  output       out2,
  output       out3,
  output       out4,
  output [7:0] out5,
  output [5:0] out6,
  output       out7
);
  assign out1 = 1'h0;
  assign out2 = 1'h0;
  assign out3 = 1'h0;
  assign out4 = 1'h1;
  assign out5 = 1'h0;
  assign out6 = 1'h0;
  assign out7 = 1'h0;
endmodule
