module Casting (
  output signed [2:0] out0,
  output        [2:0] out1,
  output        [2:0] out2
);
  assign out0 = -3'sh1;
  assign out1 = 3'h7;
  assign out2 = 3'h1;
endmodule
