module ArrayVecCase (
  input  [6:0] x_in[0:3][0:7],
  output [6:0] x_out[0:3][0:7],
  input  [5:0] y_in[0:1][0:3],
  output [5:0] y_out[0:1][0:3]
);
  ArrayVecSub u_sub (
    .x_in_0_0  ( x_in[0][0]  ),
    .x_in_0_1  ( x_in[0][1]  ),
    .x_in_0_2  ( x_in[0][2]  ),
    .x_in_0_3  ( x_in[0][3]  ),
    .x_in_0_4  ( x_in[0][4]  ),
    .x_in_0_5  ( x_in[0][5]  ),
    .x_in_0_6  ( x_in[0][6]  ),
    .x_in_0_7  ( x_in[0][7]  ),
    .x_in_1_0  ( x_in[1][0]  ),
    .x_in_1_1  ( x_in[1][1]  ),
    .x_in_1_2  ( x_in[1][2]  ),
    .x_in_1_3  ( x_in[1][3]  ),
    .x_in_1_4  ( x_in[1][4]  ),
    .x_in_1_5  ( x_in[1][5]  ),
    .x_in_1_6  ( x_in[1][6]  ),
    .x_in_1_7  ( x_in[1][7]  ),
    .x_in_2_0  ( x_in[2][0]  ),
    .x_in_2_1  ( x_in[2][1]  ),
    .x_in_2_2  ( x_in[2][2]  ),
    .x_in_2_3  ( x_in[2][3]  ),
    .x_in_2_4  ( x_in[2][4]  ),
    .x_in_2_5  ( x_in[2][5]  ),
    .x_in_2_6  ( x_in[2][6]  ),
    .x_in_2_7  ( x_in[2][7]  ),
    .x_in_3_0  ( x_in[3][0]  ),
    .x_in_3_1  ( x_in[3][1]  ),
    .x_in_3_2  ( x_in[3][2]  ),
    .x_in_3_3  ( x_in[3][3]  ),
    .x_in_3_4  ( x_in[3][4]  ),
    .x_in_3_5  ( x_in[3][5]  ),
    .x_in_3_6  ( x_in[3][6]  ),
    .x_in_3_7  ( x_in[3][7]  ),
    .x_out_0_0 ( x_out[0][0] ),
    .x_out_0_1 ( x_out[0][1] ),
    .x_out_0_2 ( x_out[0][2] ),
    .x_out_0_3 ( x_out[0][3] ),
    .x_out_0_4 ( x_out[0][4] ),
    .x_out_0_5 ( x_out[0][5] ),
    .x_out_0_6 ( x_out[0][6] ),
    .x_out_0_7 ( x_out[0][7] ),
    .x_out_1_0 ( x_out[1][0] ),
    .x_out_1_1 ( x_out[1][1] ),
    .x_out_1_2 ( x_out[1][2] ),
    .x_out_1_3 ( x_out[1][3] ),
    .x_out_1_4 ( x_out[1][4] ),
    .x_out_1_5 ( x_out[1][5] ),
    .x_out_1_6 ( x_out[1][6] ),
    .x_out_1_7 ( x_out[1][7] ),
    .x_out_2_0 ( x_out[2][0] ),
    .x_out_2_1 ( x_out[2][1] ),
    .x_out_2_2 ( x_out[2][2] ),
    .x_out_2_3 ( x_out[2][3] ),
    .x_out_2_4 ( x_out[2][4] ),
    .x_out_2_5 ( x_out[2][5] ),
    .x_out_2_6 ( x_out[2][6] ),
    .x_out_2_7 ( x_out[2][7] ),
    .x_out_3_0 ( x_out[3][0] ),
    .x_out_3_1 ( x_out[3][1] ),
    .x_out_3_2 ( x_out[3][2] ),
    .x_out_3_3 ( x_out[3][3] ),
    .x_out_3_4 ( x_out[3][4] ),
    .x_out_3_5 ( x_out[3][5] ),
    .x_out_3_6 ( x_out[3][6] ),
    .x_out_3_7 ( x_out[3][7] ),
    .y_in_0_0  ( y_in[0][0]  ),
    .y_in_0_1  ( y_in[0][1]  ),
    .y_in_0_2  ( y_in[0][2]  ),
    .y_in_0_3  ( y_in[0][3]  ),
    .y_in_1_0  ( y_in[1][0]  ),
    .y_in_1_1  ( y_in[1][1]  ),
    .y_in_1_2  ( y_in[1][2]  ),
    .y_in_1_3  ( y_in[1][3]  ),
    .y_out_0_0 ( y_out[0][0] ),
    .y_out_0_1 ( y_out[0][1] ),
    .y_out_0_2 ( y_out[0][2] ),
    .y_out_0_3 ( y_out[0][3] ),
    .y_out_1_0 ( y_out[1][0] ),
    .y_out_1_1 ( y_out[1][1] ),
    .y_out_1_2 ( y_out[1][2] ),
    .y_out_1_3 ( y_out[1][3] )
  );
endmodule
