module VecBundleCase (
  input  [15:0] io_inPacket_tx_header_0,
  input  [15:0] io_inPacket_tx_addr_0,
  input  [31:0] io_inPacket_tx_data_0,
  input  [15:0] io_inPacket_tx_header_1,
  input  [15:0] io_inPacket_tx_addr_1,
  input  [31:0] io_inPacket_tx_data_1,
  input  [15:0] io_inPacket_tx_header_2,
  input  [15:0] io_inPacket_tx_addr_2,
  input  [31:0] io_inPacket_tx_data_2,
  output [15:0] io_outPacket_rx_header_0,
  output [15:0] io_outPacket_rx_addr_0,
  output [31:0] io_outPacket_rx_data_0,
  output [15:0] io_outPacket_rx_header_1,
  output [15:0] io_outPacket_rx_addr_1,
  output [31:0] io_outPacket_rx_data_1,
  output [15:0] io_outPacket_rx_header_2,
  output [15:0] io_outPacket_rx_addr_2,
  output [31:0] io_outPacket_rx_data_2,
  output [15:0] io_outPacket_rx_header_3,
  output [15:0] io_outPacket_rx_addr_3,
  output [31:0] io_outPacket_rx_data_3
);
endmodule
