module BooleanType (
  output out0,
  output out1,
  output out2,
  output out3
);
  assign out0 = 1'h1;
  assign out1 = 1'h0;
  assign out2 = 1'h1;
  assign out3 = 1'h0;
endmodule
